//==============================================================================
// VESA Timing Generator Testbench
// 
// 自动生成时间: 2025-12-17 09:39:56
// 生成工具: VESA 视频时序计算器
//==============================================================================

`timescale 1ns / 1ps

module tb_vesa_timing_2560x1440_60hz;

//==============================================================================
// 参数定义
//==============================================================================

localparam CLK_PERIOD = 3.922;  // 时钟周期 (ns)
localparam H_TOTAL = 2848;
localparam V_TOTAL = 1492;

//==============================================================================
// 信号声明
//==============================================================================

reg         clk;
reg         rst_n;

wire        hsync;
wire        vsync;
wire        de;
wire        frame_valid;
wire [15:0] h_count;
wire [15:0] v_count;

//==============================================================================
// 时钟生成
//==============================================================================

initial begin
    clk = 1'b0;
    forever #(CLK_PERIOD/2) clk = ~clk;
end

//==============================================================================
// 复位生成
//==============================================================================

initial begin
    rst_n = 1'b0;
    #(CLK_PERIOD * 10);
    rst_n = 1'b1;
end

//==============================================================================
// 实例化被测模块
//==============================================================================

vesa_timing_2560x1440_60hz u_vesa_timing_2560x1440_60hz (
    .clk         (clk),
    .rst_n       (rst_n),
    .hsync       (hsync),
    .vsync       (vsync),
    .de          (de),
    .frame_valid (frame_valid),
    .h_count     (h_count),
    .v_count     (v_count)
);

//==============================================================================
// 监控和显示
//==============================================================================

integer frame_count;

initial begin
    frame_count = 0;
    
    // 等待复位完成
    @(posedge rst_n);
    
    // 监控帧同步信号
    forever begin
        @(negedge vsync);
        frame_count = frame_count + 1;
        $display("Time: %t ns - Frame %0d started", $time, frame_count);
        
        // 模拟 3 帧后停止
        if (frame_count >= 3) begin
            #(CLK_PERIOD * H_TOTAL * 10);
            $display("\nSimulation completed successfully!");
            $display("Total frames simulated: %0d", frame_count);
            $finish;
        end
    end
end

//==============================================================================
// 波形转储 (可选)
//==============================================================================

initial begin
    $dumpfile("tb_vesa_timing_2560x1440_60hz.vcd");
    $dumpvars(0, tb_vesa_timing_2560x1440_60hz);
end

//==============================================================================
// 超时保护
//==============================================================================

initial begin
    #(CLK_PERIOD * H_TOTAL * V_TOTAL * 5);  // 5 帧的时间
    $display("ERROR: Simulation timeout!");
    $finish;
end

endmodule
